// nios.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios (
		input  wire        clk_clk,                              //                           clk.clk
		output wire [7:0]  recv_addr_external_connection_export, // recv_addr_external_connection.export
		input  wire [31:0] recv_data_external_connection_export, // recv_data_external_connection.export
		output wire [7:0]  send_addr_external_connection_export, // send_addr_external_connection.export
		output wire [31:0] send_data_external_connection_export, // send_data_external_connection.export
		output wire [27:0] seven_seg_external_connection_export  // seven_seg_external_connection.export
	);

	wire         nios2_gen2_0_debug_reset_request_reset;                     // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [13:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                     // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [13:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;              // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;           // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;             // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;              // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;           // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;            // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_recv_data_s1_readdata;                    // recv_data:readdata -> mm_interconnect_0:recv_data_s1_readdata
	wire   [1:0] mm_interconnect_0_recv_data_s1_address;                     // mm_interconnect_0:recv_data_s1_address -> recv_data:address
	wire         mm_interconnect_0_send_addr_s1_chipselect;                  // mm_interconnect_0:send_addr_s1_chipselect -> send_addr:chipselect
	wire  [31:0] mm_interconnect_0_send_addr_s1_readdata;                    // send_addr:readdata -> mm_interconnect_0:send_addr_s1_readdata
	wire   [1:0] mm_interconnect_0_send_addr_s1_address;                     // mm_interconnect_0:send_addr_s1_address -> send_addr:address
	wire         mm_interconnect_0_send_addr_s1_write;                       // mm_interconnect_0:send_addr_s1_write -> send_addr:write_n
	wire  [31:0] mm_interconnect_0_send_addr_s1_writedata;                   // mm_interconnect_0:send_addr_s1_writedata -> send_addr:writedata
	wire         mm_interconnect_0_recv_addr_s1_chipselect;                  // mm_interconnect_0:recv_addr_s1_chipselect -> recv_addr:chipselect
	wire  [31:0] mm_interconnect_0_recv_addr_s1_readdata;                    // recv_addr:readdata -> mm_interconnect_0:recv_addr_s1_readdata
	wire   [1:0] mm_interconnect_0_recv_addr_s1_address;                     // mm_interconnect_0:recv_addr_s1_address -> recv_addr:address
	wire         mm_interconnect_0_recv_addr_s1_write;                       // mm_interconnect_0:recv_addr_s1_write -> recv_addr:write_n
	wire  [31:0] mm_interconnect_0_recv_addr_s1_writedata;                   // mm_interconnect_0:recv_addr_s1_writedata -> recv_addr:writedata
	wire         mm_interconnect_0_send_data_s1_chipselect;                  // mm_interconnect_0:send_data_s1_chipselect -> send_data:chipselect
	wire  [31:0] mm_interconnect_0_send_data_s1_readdata;                    // send_data:readdata -> mm_interconnect_0:send_data_s1_readdata
	wire   [1:0] mm_interconnect_0_send_data_s1_address;                     // mm_interconnect_0:send_data_s1_address -> send_data:address
	wire         mm_interconnect_0_send_data_s1_write;                       // mm_interconnect_0:send_data_s1_write -> send_data:write_n
	wire  [31:0] mm_interconnect_0_send_data_s1_writedata;                   // mm_interconnect_0:send_data_s1_writedata -> send_data:writedata
	wire         mm_interconnect_0_seven_seg_s1_chipselect;                  // mm_interconnect_0:seven_seg_s1_chipselect -> seven_seg:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_s1_readdata;                    // seven_seg:readdata -> mm_interconnect_0:seven_seg_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_s1_address;                     // mm_interconnect_0:seven_seg_s1_address -> seven_seg:address
	wire         mm_interconnect_0_seven_seg_s1_write;                       // mm_interconnect_0:seven_seg_s1_write -> seven_seg:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_s1_writedata;                   // mm_interconnect_0:seven_seg_s1_writedata -> seven_seg:writedata
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [mm_interconnect_0:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, onchip_memory2_0:reset, recv_addr:reset_n, recv_data:reset_n, rst_translator_001:in_reset, send_addr:reset_n, send_data:reset_n, seven_seg:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                     // rst_controller_001:reset_req -> [onchip_memory2_0:reset_req, rst_translator_001:reset_req_in]

	nios_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios_recv_addr recv_addr (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_recv_addr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_recv_addr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_recv_addr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_recv_addr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_recv_addr_s1_readdata),   //                    .readdata
		.out_port   (recv_addr_external_connection_export)       // external_connection.export
	);

	nios_recv_data recv_data (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_recv_data_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_recv_data_s1_readdata), //                    .readdata
		.in_port  (recv_data_external_connection_export)     // external_connection.export
	);

	nios_recv_addr send_addr (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_send_addr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_send_addr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_send_addr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_send_addr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_send_addr_s1_readdata),   //                    .readdata
		.out_port   (send_addr_external_connection_export)       // external_connection.export
	);

	nios_send_data send_data (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_send_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_send_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_send_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_send_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_send_data_s1_readdata),   //                    .readdata
		.out_port   (send_data_external_connection_export)       // external_connection.export
	);

	nios_seven_seg seven_seg (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_external_connection_export)       // external_connection.export
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                       (clk_clk),                                                    //                                     clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                             //      nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                         // onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                    (nios2_gen2_0_data_master_address),                           //                      nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                (nios2_gen2_0_data_master_waitrequest),                       //                                              .waitrequest
		.nios2_gen2_0_data_master_byteenable                 (nios2_gen2_0_data_master_byteenable),                        //                                              .byteenable
		.nios2_gen2_0_data_master_read                       (nios2_gen2_0_data_master_read),                              //                                              .read
		.nios2_gen2_0_data_master_readdata                   (nios2_gen2_0_data_master_readdata),                          //                                              .readdata
		.nios2_gen2_0_data_master_readdatavalid              (nios2_gen2_0_data_master_readdatavalid),                     //                                              .readdatavalid
		.nios2_gen2_0_data_master_write                      (nios2_gen2_0_data_master_write),                             //                                              .write
		.nios2_gen2_0_data_master_writedata                  (nios2_gen2_0_data_master_writedata),                         //                                              .writedata
		.nios2_gen2_0_data_master_debugaccess                (nios2_gen2_0_data_master_debugaccess),                       //                                              .debugaccess
		.nios2_gen2_0_instruction_master_address             (nios2_gen2_0_instruction_master_address),                    //               nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest         (nios2_gen2_0_instruction_master_waitrequest),                //                                              .waitrequest
		.nios2_gen2_0_instruction_master_read                (nios2_gen2_0_instruction_master_read),                       //                                              .read
		.nios2_gen2_0_instruction_master_readdata            (nios2_gen2_0_instruction_master_readdata),                   //                                              .readdata
		.nios2_gen2_0_instruction_master_readdatavalid       (nios2_gen2_0_instruction_master_readdatavalid),              //                                              .readdatavalid
		.nios2_gen2_0_debug_mem_slave_address                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //                  nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                              .write
		.nios2_gen2_0_debug_mem_slave_read                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                              .read
		.nios2_gen2_0_debug_mem_slave_readdata               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                              .readdata
		.nios2_gen2_0_debug_mem_slave_writedata              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                              .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                              .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                              .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                              .debugaccess
		.onchip_memory2_0_s1_address                         (mm_interconnect_0_onchip_memory2_0_s1_address),              //                           onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                           (mm_interconnect_0_onchip_memory2_0_s1_write),                //                                              .write
		.onchip_memory2_0_s1_readdata                        (mm_interconnect_0_onchip_memory2_0_s1_readdata),             //                                              .readdata
		.onchip_memory2_0_s1_writedata                       (mm_interconnect_0_onchip_memory2_0_s1_writedata),            //                                              .writedata
		.onchip_memory2_0_s1_byteenable                      (mm_interconnect_0_onchip_memory2_0_s1_byteenable),           //                                              .byteenable
		.onchip_memory2_0_s1_chipselect                      (mm_interconnect_0_onchip_memory2_0_s1_chipselect),           //                                              .chipselect
		.onchip_memory2_0_s1_clken                           (mm_interconnect_0_onchip_memory2_0_s1_clken),                //                                              .clken
		.recv_addr_s1_address                                (mm_interconnect_0_recv_addr_s1_address),                     //                                  recv_addr_s1.address
		.recv_addr_s1_write                                  (mm_interconnect_0_recv_addr_s1_write),                       //                                              .write
		.recv_addr_s1_readdata                               (mm_interconnect_0_recv_addr_s1_readdata),                    //                                              .readdata
		.recv_addr_s1_writedata                              (mm_interconnect_0_recv_addr_s1_writedata),                   //                                              .writedata
		.recv_addr_s1_chipselect                             (mm_interconnect_0_recv_addr_s1_chipselect),                  //                                              .chipselect
		.recv_data_s1_address                                (mm_interconnect_0_recv_data_s1_address),                     //                                  recv_data_s1.address
		.recv_data_s1_readdata                               (mm_interconnect_0_recv_data_s1_readdata),                    //                                              .readdata
		.send_addr_s1_address                                (mm_interconnect_0_send_addr_s1_address),                     //                                  send_addr_s1.address
		.send_addr_s1_write                                  (mm_interconnect_0_send_addr_s1_write),                       //                                              .write
		.send_addr_s1_readdata                               (mm_interconnect_0_send_addr_s1_readdata),                    //                                              .readdata
		.send_addr_s1_writedata                              (mm_interconnect_0_send_addr_s1_writedata),                   //                                              .writedata
		.send_addr_s1_chipselect                             (mm_interconnect_0_send_addr_s1_chipselect),                  //                                              .chipselect
		.send_data_s1_address                                (mm_interconnect_0_send_data_s1_address),                     //                                  send_data_s1.address
		.send_data_s1_write                                  (mm_interconnect_0_send_data_s1_write),                       //                                              .write
		.send_data_s1_readdata                               (mm_interconnect_0_send_data_s1_readdata),                    //                                              .readdata
		.send_data_s1_writedata                              (mm_interconnect_0_send_data_s1_writedata),                   //                                              .writedata
		.send_data_s1_chipselect                             (mm_interconnect_0_send_data_s1_chipselect),                  //                                              .chipselect
		.seven_seg_s1_address                                (mm_interconnect_0_seven_seg_s1_address),                     //                                  seven_seg_s1.address
		.seven_seg_s1_write                                  (mm_interconnect_0_seven_seg_s1_write),                       //                                              .write
		.seven_seg_s1_readdata                               (mm_interconnect_0_seven_seg_s1_readdata),                    //                                              .readdata
		.seven_seg_s1_writedata                              (mm_interconnect_0_seven_seg_s1_writedata),                   //                                              .writedata
		.seven_seg_s1_chipselect                             (mm_interconnect_0_seven_seg_s1_chipselect)                   //                                              .chipselect
	);

	nios_irq_mapper irq_mapper (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
