-- megafunction wizard: %RAM: 1-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: DM_RAM.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Standard Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY DM_RAM IS
	PORT
	(
		address		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
		clock		: IN STD_LOGIC  := '1';
		data		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		wren		: IN STD_LOGIC ;
		q		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END DM_RAM;


ARCHITECTURE SYN OF dm_ram IS
	type slv_array_t is array (natural range <>) of std_logic_vector(15 downto 0);

	signal mux_signals : slv_array_t(0 to 15);
	signal sel_z_internal : integer;
	signal write_z : std_logic_vector(0 to 15);
	signal sel_z : std_logic_vector(3 downto 0);

BEGIN
	REG_FILE :
	for I in 0 to 15 generate
		REGX : entity work.REG1_GENERIC
		generic map(
			LEN => 16
		)
		port map(
			reg_in => data, 
			writ => write_z(i),
			reset => '0',
			clk => clock,
			reg_out => mux_signals(i)
		);
	end generate REG_FILE;

	sel_z <= address(3 downto 0);

    process(sel_z, wren)
    begin
        write_z <= (others => '0');
        write_z(to_integer(unsigned(sel_z))) <= wren;
    end process;

    q <= mux_signals(to_integer(unsigned(sel_z)));

END SYN;
